package Soc where

import Utils
import GetPut
import ClientServer
import Connectable

import Vector
import AXI4
import AXI4_Lite
import AXI4_Lite_Adapter

import TestBench
import UART

import Core
import CoreOOO
import Screen
import SdCard
import Clint

--import CC
import LSU
import BCache
import BranchPred
import SDRAM

interface CPU_IFC =
  memory :: PinsSDRAM {-# prefix="" #-}
  led :: Bit 8 {-# always_ready, always_enabled #-}
  ftdi_rxd :: Bit 1 {-# always_ready, always_enabled #-}
  ftdi_txd :: Bit 1 -> Action {-# always_ready, always_enabled, arg_names= [ftdi_txd], prefix="" #-}
  vga_out :: VGAFabric {-# prefix = "" #-}
  btn_in :: Bit 6 -> Action {-# always_ready, always_enabled, arg_names= [btn], prefix = "" #-}
  sdcard_fab :: SdCardFab {-# prefix = "sd" #-}

{-# verilog mkCPU #-}
mkCPU :: Module CPU_IFC
mkCPU = module
  sdram <- mkSdramAXI4 32'h80000000
  let wr_port = sdram.slave.write
  let rd_port = sdram.slave.read
  -- wr_port <- mkWrAXI4_Master Pipeline
  -- rd_port <- mkRdAXI4_Master Pipeline

  core <- mkCoreOOO
  let core_i_rd = core.rd_imem

  let alloc_size :: Integer = 0x3d6f -- 32'h800 -- 32'h660 -- 32'h23000
  let offset :: Bit 32 = 32'h80000000
  let is_vga :: Bit 32 -> Bool = \x -> x >= 32'h40000000 && x < 32'h50000000
  let is_btn :: Bit 32 -> Bool = \x -> x == 32'h20000000
  let is_sdcard :: Bit 32 -> Bool = \x -> x == 32'h50000000
  let is_clint :: Bit 32 -> Bool = \x -> x >= 32'h30000000 && x < 32'h3000C000

  rom <- mkRom (RomConfig{name="Mem.hex"; start=offset; size=alloc_size; maxPhase=0})
  clint <- mkCLINT_AXI4_Lite 32'h30000000
  vga <- mkVGA_AXI4_Lite 32'h40000000
  sdcard <- mkSdCard 32'h50000000
  uart <- mkUART 217 32'h10000000
  btn <- mkBtn 32'h20000000

  let rd_masters_lite :: Vector 1 (RdAXI4_Lite_Master 32 4) = core.rd_mmio :> nil
  let wr_masters_lite :: Vector 1 (WrAXI4_Lite_Master 32 4) = core.wr_mmio :> nil

  let rd_slaves_lite :: Vector 5 (RdAXI4_Lite_Slave 32 4) =
        uart.axi4.read :> vga.axi4.read :> btn.axi4.read
        :> clint.read :> sdcard.axi4.read :> nil
  let wr_slaves_lite :: Vector 5 (WrAXI4_Lite_Slave 32 4) =
        uart.axi4.write :> vga.axi4.write :> btn.axi4.write
        :> clint.write :> sdcard.axi4.write :> nil

  let rdReqLiteDispatch :: AXI4_Lite_RRequest 32 -> Bit 3 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_vga req.addr then 1 else
        if is_btn req.addr then 2 else
        if is_clint req.addr then 3 else
        if is_sdcard req.addr then 4 else 0
  let wrReqLiteDispatch :: AXI4_Lite_WRequest 32 4 -> Bit 3 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_vga req.addr then 1 else
        if is_btn req.addr then 2 else
        if is_clint req.addr then 3 else
        if is_sdcard req.addr then 4 else 0

  mkXBarRdAXI4_Lite rd_masters_lite rd_slaves_lite rdReqLiteDispatch
  mkXBarWrAXI4_Lite wr_masters_lite wr_slaves_lite wrReqLiteDispatch

  let rd_masters :: Vector 2 (RdAXI4_Master 4 32 4) = core.rd_dmem :> core_i_rd :> nil
  let wr_masters :: Vector 1 (WrAXI4_Master 4 32 4) = core.wr_dmem :> nil

  let rd_slaves :: Vector 2 (RdAXI4_Slave 4 32 4) = rom.read :> rd_port :> nil
  let wr_slaves :: Vector 2 (WrAXI4_Slave 4 32 4) = rom.write :> wr_port :> nil

  let rdReqDispatch :: AXI4_RRequest 4 32 -> Bit 1 =
        \ req -> if req.addr < offset || req.addr >= offset + fromInteger alloc_size then 1 else 0
  let wrReqDispatch :: AXI4_AWRequest 4 32 -> Bit 1 =
        \ req -> if req.addr < offset || req.addr >= offset + fromInteger alloc_size then 1 else 0

  mkXBarRdAXI4 rd_masters rd_slaves rdReqDispatch
  mkXBarWrAXI4 wr_masters wr_slaves wrReqDispatch

  rules
    "uart interrupt": when True ==> do
      core.set_meip(True)
      uart.interrupt

    "btn interrupt": when True ==> do
      core.set_meip(True)
      btn.interrupt

    "clint timer interrupt": when True ==> do
      core.set_mtip(clint.timer_interrupt)

    "clint software interrupt": when True ==> do
      core.set_msip(clint.software_interrupt)

  interface
    memory = sdram.memory
    sdcard_fab = sdcard.fabric
    ftdi_rxd = uart.transmit
    ftdi_txd = uart.receive
    vga_out = vga.fabric
    btn_in = btn.fabric
    led = uart.leds

{-# verilog mkCPU #-}
mkCPU_SIM :: Module Empty
mkCPU_SIM = module
  sdram <- mkSdramAXI4 32'h80000000
  let wr_port = sdram.slave.write
  let rd_port = sdram.slave.read

  core <- mkCoreOOO
  let core_i_rd = core.rd_imem

  let alloc_size :: Integer = 300000 --33 * 1024 * 1024 -- maxBound
  let offset :: Bit 32 = 32'h80000000
  let is_vga :: Bit 32 -> Bool = \x -> x >= 32'h40000000 && x < 32'h50000000
  let is_btn :: Bit 32 -> Bool = \x -> x == 32'h20000000
  let is_clint :: Bit 32 -> Bool = \x -> x >= 32'h30000000 && x < 32'h3000C000
  let is_sdcard :: Bit 32 -> Bool = \x -> x == 32'h50000000

  rom <- mkRom (RomConfig{name="Mem.hex"; start=offset; size=alloc_size; maxPhase=0})
  clint <- mkCLINT_AXI4_Lite 32'h30000000
  vga <- mkVGA_AXI4_Lite 32'h40000000
  sdcard <- mkSdCard 32'h50000000
  uart <- mkUART 217 32'h10000000
  btn <- mkBtn 32'h20000000

  let rd_masters_lite :: Vector 1 (RdAXI4_Lite_Master 32 4) = core.rd_mmio :> nil
  let wr_masters_lite :: Vector 1 (WrAXI4_Lite_Master 32 4) = core.wr_mmio :> nil

  let rd_slaves_lite :: Vector 5 (RdAXI4_Lite_Slave 32 4) =
        uart.axi4.read :> vga.axi4.read :> btn.axi4.read
        :> clint.read :> sdcard.axi4.read :> nil
  let wr_slaves_lite :: Vector 5 (WrAXI4_Lite_Slave 32 4) =
        uart.axi4.write :> vga.axi4.write :> btn.axi4.write
        :> clint.write :> sdcard.axi4.write :> nil

  let rdReqLiteDispatch :: AXI4_Lite_RRequest 32 -> Bit 3 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_vga req.addr then 1 else
        if is_clint req.addr then 3 else
        if is_btn req.addr then 2 else
        if is_sdcard req.addr then 4 else 0
  let wrReqLiteDispatch :: AXI4_Lite_WRequest 32 4 -> Bit 3 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_vga req.addr then 1 else
        if is_clint req.addr then 3 else
        if is_btn req.addr then 2 else
        if is_sdcard req.addr then 4 else 0

  mkXBarRdAXI4_Lite rd_masters_lite rd_slaves_lite rdReqLiteDispatch
  mkXBarWrAXI4_Lite wr_masters_lite wr_slaves_lite wrReqLiteDispatch

  let rd_masters :: Vector 2 (RdAXI4_Master 4 32 4) = core.rd_dmem :> core_i_rd :> nil
  let wr_masters :: Vector 1 (WrAXI4_Master 4 32 4) = core.wr_dmem :> nil

  let rd_slaves :: Vector 2 (RdAXI4_Slave 4 32 4) = rom.read :> rd_port :> nil
  let wr_slaves :: Vector 2 (WrAXI4_Slave 4 32 4) = rom.write :> wr_port :> nil

  let rdReqDispatch :: AXI4_RRequest 4 32 -> Bit 1 =
        \ req -> if req.addr < offset || req.addr >= offset + fromInteger alloc_size then 1 else 0
  let wrReqDispatch :: AXI4_AWRequest 4 32 -> Bit 1 =
        \ req -> if req.addr < offset || req.addr >= offset + fromInteger alloc_size then 1 else 0

  mkXBarRdAXI4 rd_masters rd_slaves rdReqDispatch
  mkXBarWrAXI4 wr_masters wr_slaves wrReqDispatch

  cycle :: Reg (Bit 32) <- mkReg 0

  rules
    "give sdram data": when True ==> do
      sdram.memory.sdram_d_in 0

    "cycle count": when True ==> do
      cycle := cycle + 1

    "uart interrupt": when False ==> do
      core.set_meip(True)
      uart.interrupt

    "btn interrupt": when False ==> do
      core.set_meip(True)
      --btn.interrupt

    "receive_uart": when True ==> do
      uart.receive 1

    "receive btn": when True ==> do
      btn.fabric 0

    "sdcard receive": when True ==> do
      sdcard.fabric.cmd_in 0
      sdcard.fabric.data_in 0

    "clint timer interrupt": when True ==> do
      core.set_mtip(clint.timer_interrupt)

    "clint software interrupt": when True ==> do
      core.set_msip(clint.software_interrupt)

interface CPU_MINIMAL_IFC =
  led :: Bit 8 {-# always_ready, always_enabled #-}
  ftdi_rxd :: Bit 1 {-# always_ready, always_enabled #-}
  ftdi_txd :: Bit 1 -> Action {-# always_ready, always_enabled, arg_names= [ftdi_txd], prefix="" #-}
  -- write SDRAM port using AXI4 protocol
  wr_axi4 :: WrAXI4_Master_Fab 4 32 4 {-# prefix="" #-}
  -- read SDRAM port using AXI4 protocol
  rd_axi4 :: RdAXI4_Master_Fab 4 32 4 {-# prefix="" #-}

{-# verilog mkCPU #-}
mkCPU_MINIMAL :: Module CPU_MINIMAL_IFC
mkCPU_MINIMAL = module
  wr_port <- mkWrAXI4_Master Pipeline
  rd_port <- mkRdAXI4_Master Pipeline

  core <- mkCoreOOO
  let core_i_rd = core.rd_imem

  let alloc_size :: Integer = 0x3d6f -- 32'h800 -- 32'h660 -- 32'h23000
  let offset :: Bit 32 = 32'h80000000
  let is_clint :: Bit 32 -> Bool = \x -> x >= 32'h30000000 && x < 32'h3000C000

  rom <- mkRom (RomConfig{name="Mem.mem"; start=offset; size=alloc_size; maxPhase=0})
  clint <- mkCLINT_AXI4_Lite 32'h30000000
  uart <- mkUART 347 32'h10000000

  let rd_masters_lite :: Vector 1 (RdAXI4_Lite_Master 32 4) = core.rd_mmio :> nil
  let wr_masters_lite :: Vector 1 (WrAXI4_Lite_Master 32 4) = core.wr_mmio :> nil

  let rd_slaves_lite :: Vector 2 (RdAXI4_Lite_Slave 32 4) =
        uart.axi4.read :> clint.read :> nil
  let wr_slaves_lite :: Vector 2 (WrAXI4_Lite_Slave 32 4) =
        uart.axi4.write :> clint.write :> nil

  let rdReqLiteDispatch :: AXI4_Lite_RRequest 32 -> Bit 1 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_clint req.addr then 1 else 0
  let wrReqLiteDispatch :: AXI4_Lite_WRequest 32 4 -> Bit 1 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_clint req.addr then 1 else 0

  mkXBarRdAXI4_Lite rd_masters_lite rd_slaves_lite rdReqLiteDispatch
  mkXBarWrAXI4_Lite wr_masters_lite wr_slaves_lite wrReqLiteDispatch

  let rd_masters :: Vector 2 (RdAXI4_Master 4 32 4) = core.rd_dmem :> core_i_rd :> nil
  let wr_masters :: Vector 1 (WrAXI4_Master 4 32 4) = core.wr_dmem :> nil

  let rd_slaves :: Vector 2 (RdAXI4_Slave 4 32 4) = rom.read :> rd_port.server :> nil
  let wr_slaves :: Vector 2 (WrAXI4_Slave 4 32 4) = rom.write :> wr_port.server :> nil

  let rdReqDispatch :: AXI4_RRequest 4 32 -> Bit 1 =
        \ req -> if req.addr < offset || req.addr >= offset + fromInteger alloc_size then 1 else 0
  let wrReqDispatch :: AXI4_AWRequest 4 32 -> Bit 1 =
        \ req -> if req.addr < offset || req.addr >= offset + fromInteger alloc_size then 1 else 0

  mkXBarRdAXI4 rd_masters rd_slaves rdReqDispatch
  mkXBarWrAXI4 wr_masters wr_slaves wrReqDispatch

  rules
    "uart interrupt": when True ==> do
      core.set_meip(True)
      uart.interrupt

    "clint timer interrupt": when True ==> do
      core.set_mtip(clint.timer_interrupt)

    "clint software interrupt": when True ==> do
      core.set_msip(clint.software_interrupt)

  interface
    wr_axi4 = wr_port.fabric
    rd_axi4 = rd_port.fabric
    ftdi_rxd = uart.transmit
    ftdi_txd = uart.receive
    led = uart.leds


interface CPU_NO_SDRAM_IFC =
  led :: Bit 8 {-# always_ready, always_enabled #-}
  ftdi_rxd :: Bit 1 {-# always_ready, always_enabled #-}
  ftdi_txd :: Bit 1 -> Action {-# always_ready, always_enabled, arg_names= [ftdi_txd], prefix="" #-}

{-# verilog mkCPU #-}
mkCPU_NO_SDRAM :: Module CPU_NO_SDRAM_IFC
mkCPU_NO_SDRAM  = module
  core <- mkCoreOOO
  let core_i_rd = core.rd_imem

  let alloc_size :: Integer = 0x3d6f -- 32'h800 -- 32'h660 -- 32'h23000
  let offset :: Bit 32 = 32'h80000000
  let is_clint :: Bit 32 -> Bool = \x -> x >= 32'h30000000 && x < 32'h3000C000

  rom <- mkRom (RomConfig{name="Mem.mem"; start=offset; size=alloc_size; maxPhase=0})
  clint <- mkCLINT_AXI4_Lite 32'h30000000
  uart <- mkUART 347 32'h10000000

  let rd_masters_lite :: Vector 1 (RdAXI4_Lite_Master 32 4) = core.rd_mmio :> nil
  let wr_masters_lite :: Vector 1 (WrAXI4_Lite_Master 32 4) = core.wr_mmio :> nil

  let rd_slaves_lite :: Vector 2 (RdAXI4_Lite_Slave 32 4) =
        uart.axi4.read :> clint.read :> nil
  let wr_slaves_lite :: Vector 2 (WrAXI4_Lite_Slave 32 4) =
        uart.axi4.write :> clint.write :> nil

  let rdReqLiteDispatch :: AXI4_Lite_RRequest 32 -> Bit 1 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_clint req.addr then 1 else 0
  let wrReqLiteDispatch :: AXI4_Lite_WRequest 32 4 -> Bit 1 =
        \ req -> if req.addr == 32'h10000000 then 0 else
        if is_clint req.addr then 1 else 0

  mkXBarRdAXI4_Lite rd_masters_lite rd_slaves_lite rdReqLiteDispatch
  mkXBarWrAXI4_Lite wr_masters_lite wr_slaves_lite wrReqLiteDispatch

  let rd_masters :: Vector 2 (RdAXI4_Master 4 32 4) = core.rd_dmem :> core_i_rd :> nil
  let wr_masters :: Vector 1 (WrAXI4_Master 4 32 4) = core.wr_dmem :> nil

  let rd_slaves :: Vector 1 (RdAXI4_Slave 4 32 4) = rom.read :> nil
  let wr_slaves :: Vector 1 (WrAXI4_Slave 4 32 4) = rom.write :> nil

  let rdReqDispatch :: AXI4_RRequest 4 32 -> Bit 0 = \ req -> 0
  let wrReqDispatch :: AXI4_AWRequest 4 32 -> Bit 0 = \ req -> 0

  mkXBarRdAXI4 rd_masters rd_slaves rdReqDispatch
  mkXBarWrAXI4 wr_masters wr_slaves wrReqDispatch

  rules
    "uart interrupt": when True ==> do
      core.set_meip(True)
      uart.interrupt

    "clint timer interrupt": when True ==> do
      core.set_mtip(clint.timer_interrupt)

    "clint software interrupt": when True ==> do
      core.set_msip(clint.software_interrupt)

  interface
    ftdi_rxd = uart.transmit
    ftdi_txd = uart.receive
    led = uart.leds


{-# verilog mkCPU #-}
mkDDR3_TEST :: Module CPU_MINIMAL_IFC
mkDDR3_TEST = module
  wr_port <- mkWrAXI4_Master (Normal(2))
  rd_port <- mkRdAXI4_Master (Normal(2))

  tx_uart <- mkTxUART (83_000_000 / 115200)
  rx_uart <- mkRxUART (83_000_000 / 115200)

  counter :: Reg (Bit 32) <- mkReg 0

  state :: Reg (Bit 2) <- mkReg 0

  rules
    "count": when True ==> do
      counter := counter + 1

    --"testRl": when True ==> do
    --  tx_uart.put ((zeroExtend counter[27:25]) | 8'h30)

    "send_ddr3 write request": when state == 0 ==> do
      wr_port.server.awrequest.put (AXI4_AWRequest{addr=0; id=0; length=0; burst=INCR})
      wr_port.server.wrequest.put (AXI4_WRequest{bytes=7; strb=15; last=True})
      state := 1

    "receive w response": when state == 1 ==> do
      resp <- wr_port.server.response.get
      state := 2

    "send_ddr3 read request": when state == 2 && counter[26:0] == 0 ==> do
      rd_port.server.request.put (AXI4_RRequest{addr=0; id=0; length=0; burst=INCR})

    "receive ddr3 response": when True ==> do
      resp <- rd_port.server.response.get
      tx_uart.put ((zeroExtend resp.bytes[2:0]) | 8'h30)

  interface
    wr_axi4 = wr_port.fabric
    rd_axi4 = rd_port.fabric
    ftdi_rxd = tx_uart.transmit
    ftdi_txd = rx_uart.receive
    led = tx_uart.leds -- counter[27:20]
