import AXI4_Lite :: *;
import AXI4 :: *;

import Utils :: *;
import Ehr :: *;
import Fifo :: *;

