import AXI4_Lite :: *;
import GetPut :: *;
import Utils :: *;
import AXI4 :: *;
import Fifo :: *;
import Ehr :: *;
