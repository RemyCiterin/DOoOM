import ForwardRegFile :: *;
import RegFile :: *;
import Utils :: *;
import Decode :: *;
import Vector :: *;
import Fifo :: *;
import Ehr :: *;
import CSR :: *;
import OOO :: *;

// first < deq < writeBack < read < enq
interface ROB;
  /* Stage 1: enqueue */
  // read an entry from the rob
  method Maybe#(ExecOutput) read1(RobIndex index);

  // read an entry from the rob
  method Maybe#(ExecOutput) read2(RobIndex index);

  // enqueue a new entry in the reorder buffer
  method ActionValue#(RobIndex) enq(RobEntry entry);

  /* Stage 2: write back */
  // write back the result of the execution of an instruction to the rob
  method Action writeBack(RobIndex index, ExecOutput result);

  /* Stage 3: dequeue */
  // return the first element of the rob before deq
  method RobEntry first;

  // return the first index of the rob before deq
  method RobIndex first_index;

  // return the result of the execution of the first item
  method Maybe#(ExecOutput) first_result;

  // dequeue an element of the rob
  method Action deq;
endinterface

(* synthesize *)
module mkROB(ROB);
  RegFile#(RobIndex, RobEntry) data <- mkRegFileFull;
  ForwardRegFile#(RobIndex, ExecOutput) results <- mkForwardRegFileFull;
  Ehr#(2, Bit#(RobSize)) resultValid <- mkEhr(0);

  Ehr#(2, RobIndex) firstP <- mkEhr(0);
  Reg#(RobIndex) nextP <- mkReg(0);

  RobIndex max_index = fromInteger(valueOf(RobSize) - 1);

  Ehr#(2, Bool) empty <- mkEhr(True);
  Ehr#(2, Bool) full <- mkEhr(False);

  // use port 1 of data, empty and full
  method ActionValue#(RobIndex) enq(RobEntry entry)
    if (!full[1]);
    actionvalue
      resultValid[1][nextP] <= 0;
      let next_nextP = (nextP == max_index ? 0 : nextP + 1);
      let index = nextP;

      data.upd(nextP, entry);
      empty[1] <= False;
      nextP <= next_nextP;

      if (next_nextP == firstP[1])
        full[1] <= True;

      return index;
    endactionvalue
  endmethod

  method RobEntry first if (!empty[0]);
    return data.sub(firstP[0]);
  endmethod

  method RobIndex first_index if (!empty[0]);
    return firstP[0];
  endmethod

  method first_result if (!empty[0]);
    return resultValid[0][firstP[0]] == 1 ?
      Valid(results.sub(firstP[0])) : Invalid;
  endmethod

  method Action deq if (!empty[0]);
    let next_firstP = (firstP[0] == max_index ? 0 : firstP[0] + 1);
    full[0] <= False;

    firstP[0] <= next_firstP;
    if (next_firstP == nextP)
      empty[0] <= True;
  endmethod

  method Maybe#(ExecOutput) read1(RobIndex index);
    return resultValid[1][index] == 1 ?
      Valid(results.forward(index)) : Invalid;
  endmethod

  method Maybe#(ExecOutput) read2(RobIndex index);
    return resultValid[1][index] == 1 ?
      Valid(results.forward(index)) : Invalid;
  endmethod

  method Action writeBack(RobIndex index, ExecOutput result);
    action
      results.upd(index, result);
      resultValid[0][index] <= 1;
    endaction
  endmethod
endmodule
